../../submodules/marga/hdl/gpa_fhdo_iface.sv