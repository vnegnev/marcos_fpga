../../submodules/flocra/hdl/flocra.sv