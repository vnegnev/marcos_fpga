../../submodules/flocra/hdl/flodecode.sv