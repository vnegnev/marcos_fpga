../../submodules/flocra/hdl/flofifo.sv