../../submodules/flocra/hdl/flobuffer.sv