../../submodules/marga/hdl/mardecode.sv