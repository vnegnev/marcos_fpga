../../submodules/flocra/hdl/ocra1_iface.sv