../../submodules/marga/hdl/marga.sv