../../submodules/marga/hdl/ocra1_iface.sv