../../submodules/marga/hdl/marfifo.sv