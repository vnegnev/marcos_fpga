../../submodules/marga/hdl/marbuffer.sv