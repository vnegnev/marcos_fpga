../../submodules/flocra/hdl/gpa_fhdo_iface.sv